uint64_t code[] = '{
64'h2800002000a3d70a, 
64'h0000000800000000, 
64'h0000000800000000, 
64'h0000000800000000, 
64'h0000000800000000, 
64'h2400401840000000, 
64'h100080080ccccccc, 
64'h0000000800000000, 
64'h0000000800000000, 
64'h0000000800000000, 
64'h0000000800000000, 
64'hc000000800000000, 
64'h0000000800000000, 
64'h0000000800000000, 
64'h0000000800000000, 
64'h0000000800000000, 
64'h0000000800000000, 
64'h0000000800000000};
